module eightbitadder(a,b,cin,s,cout);
input [7:0]a,b;
input cin;
output [7:0]s;
output cout;
wire [7:0]c;
assign cout= c[7];
fulladd a1(a[0],b[0],cin,s[0],c[0]);
fulladd a2(a[1],b[1],c[0],s[1],c[1]);
fulladd a3(a[2],b[2],c[1],s[2],c[2]);
fulladd a4(a[3],b[3],c[2],s[3],c[3]);
fulladd a5(a[4],b[4],c[3],s[4],c[4]);
fulladd a6(a[5],b[5],c[4],s[5],c[5]);
fulladd a7(a[6],b[6],c[5],s[6],c[6]);
fulladd a8(a[7],b[7],c[6],s[7],c[7]);
endmodule
module fulladd(a,b,c,sum,carry);
input a,b,c;
output sum,carry;
assign sum=a^b^c;
assign carry=(a&b)|(a&c)|(b&c);
endmodule
