module eightbitmultiplier (x,y,p);
input [7:0]x,y;
output [15:0]p;
wire [63:0]w;
wire [54:0]c;
wire [41:0]s;
and a1 (w[0],x[0],y[0]);
and a2 (w[1],x[1],y[0]);
and a3 (w[2],x[2],y[0]);
and a4 (w[3],x[3],y[0]);
and a5 (w[4],x[4],y[0]);
and a6 (w[5],x[5],y[0]);
and a7 (w[6],x[6],y[0]);
and a8 (w[7],x[7],y[0]);
and a9 (w[8],x[0],y[1]);
and a10 (w[9],x[1],y[1]);
and a11 (w[10],x[2],y[1]);
and a12 (w[11],x[3],y[1]);
and a13 (w[12],x[4],y[1]);
and a14 (w[13],x[5],y[1]);
and a15 (w[14],x[6],y[1]);
and a16 (w[15],x[7],y[1]);
and a17 (w[16],x[0],y[2]);
and a18 (w[17],x[1],y[2]);
and a19 (w[18],x[2],y[2]);
and a20 (w[19],x[3],y[2]);
21
and a21 (w[20],x[4],y[2]);
and a22 (w[21],x[5],y[2]);
and a23 (w[22],x[6],y[2]);
and a24 (w[23],x[7],y[2]);
and a25 (w[24],x[0],y[3]);
and a26 (w[25],x[1],y[3]);
and a27 (w[26],x[2],y[3]);
and a28 (w[27],x[3],y[3]);
and a29 (w[28],x[4],y[3]);
and a30 (w[29],x[5],y[3]);
and a31 (w[30],x[6],y[3]);
and a32 (w[31],x[7],y[3]);
and a33 (w[32],x[0],y[4]);
and a34 (w[33],x[1],y[4]);
and a35 (w[34],x[2],y[4]);
and a36 (w[35],x[3],y[4]);
and a37 (w[36],x[4],y[4]);
and a38 (w[37],x[5],y[4]);
and a39 (w[38],x[6],y[4]);
and a40 (w[39],x[7],y[4]);
and a41 (w[40],x[0],y[5]);
and a42 (w[41],x[1],y[5]);
and a43 (w[42],x[2],y[5]);
and a44 (w[43],x[3],y[5]);
and a45 (w[44],x[4],y[5]);
and a46 (w[45],x[5],y[5]);
and a47 (w[46],x[6],y[5]);
and a48 (w[47],x[7],y[5]);
22
and a49 (w[48],x[0],y[6]);
and a50 (w[49],x[1],y[6]);
and a51 (w[50],x[2],y[6]);
and a52 (w[51],x[3],y[6]);
and a53 (w[52],x[4],y[6]);
and a54 (w[53],x[5],y[6]);
and a55 (w[54],x[6],y[6]);
and a56 (w[55],x[7],y[6]);
and a57 (w[56],x[0],y[7]);
and a58 (w[57],x[1],y[7]);
and a59 (w[58],x[2],y[7]);
and a60 (w[59],x[3],y[7]);
and a61 (w[60],x[4],y[7]);
and a62 (w[61],x[5],y[7]);
and a63 (w[62],x[6],y[7]);
and a64 (w[63],x[7],y[7]);
assign p[0]=w[0];
halfadd ha1(w[1],w[8],p[1],c[0]);
fulladd fa1(w[2],w[9],c[0],s[0],c[1]);
fulladd fa2(w[3],w[10],c[1],s[1],c[2]);
fulladd fa3(w[4],w[11],c[2],s[2],c[3]);
fulladd fa4(w[5],w[12],c[3],s[3],c[4]);
fulladd fa5(w[6],w[13],c[4],s[4],c[5]);
fulladd fa6(w[7],w[14],c[5],s[5],c[6]);
halfadd ha2(w[15],c[6],s[6],c[7]);
halfadd ha3(s[0],w[16],p[2],c[8]);
fulladd fa7(s[1],w[17],c[8],s[7],c[9]);
fulladd fa8(s[2],w[18],c[9],s[8],c[10]);
fulladd fa9(s[3],w[19],c[10],s[9],c[11]);
23
fulladd fa10(s[4],w[20],c[11],s[10],c[12]);
fulladd fa11(s[5],w[21],c[12],s[11],c[13]);
fulladd fa12(s[6],w[22],c[13],s[12],c[14]);
fulladd fa13(c[7],w[23],c[14],s[13],c[15]);
halfadd ha4(s[7],w[24],p[3],c[16]);
fulladd fa14(s[8],w[25],c[16],s[14],c[17]);
fulladd fa15(s[9],w[26],c[17],s[15],c[18]);
fulladd fa16(s[10],w[27],c[18],s[16],c[19]);
fulladd fa17(s[11],w[28],c[19],s[17],c[20]);
fulladd fa18(s[12],w[29],c[20],s[18],c[21]);
fulladd fa19(s[13],w[30],c[21],s[19],c[22]);
fulladd fa20(c[15],w[31],c[22],s[20],c[23]);
halfadd ha5(s[14],w[32],p[4],c[24]);
fulladd fa21(s[15],w[33],c[24],s[21],c[25]);
fulladd fa22(s[16],w[34],c[25],s[22],c[26]);
fulladd fa23(s[17],w[35],c[26],s[23],c[27]);
fulladd fa24(s[18],w[36],c[27],s[24],c[28]);
fulladd fa25(s[19],w[37],c[28],s[25],c[29]);
fulladd fa26(s[20],w[38],c[29],s[26],c[30]);
fulladd fa27(c[23],w[39],c[30],s[27],c[31]);
halfadd ha6(s[21],w[40],p[5],c[32]);
fulladd fa28(s[22],w[41],c[32],s[28],c[33]);
fulladd fa29(s[23],w[42],c[33],s[29],c[34]);
fulladd fa30(s[24],w[43],c[34],s[30],c[35]);
fulladd fa31(s[25],w[44],c[35],s[31],c[36]);
fulladd fa32(s[26],w[45],c[36],s[32],c[37]);
fulladd fa33(s[27],w[46],c[37],s[33],c[38]);
fulladd fa34(c[31],w[47],c[38],s[34],c[39]);
24
halfadd ha7(s[28],w[48],p[6],c[40]);
fulladd fa35(s[29],w[49],c[40],s[35],c[41]);
fulladd fa36(s[30],w[50],c[41],s[36],c[42]);
fulladd fa37(s[31],w[51],c[42],s[37],c[43]);
fulladd fa38(s[32],w[52],c[43],s[38],c[44]);
fulladd fa39(s[33],w[53],c[44],s[39],c[45]);
fulladd fa40(s[34],w[54],c[45],s[40],c[46]);
fulladd fa41(c[39],w[55],c[46],s[41],c[47]);
halfadd ha8(s[35],w[56],p[7],c[48]);
fulladd fa42(s[36],w[57],c[48],p[8],c[49]);
fulladd fa43(s[37],w[58],c[49],p[9],c[50]);
fulladd fa44(s[38],w[59],c[50],p[10],c[51]);
fulladd fa45(s[39],w[60],c[51],p[11],c[52]);
fulladd fa46(s[40],w[61],c[52],p[12],c[53]);
fulladd fa47(s[41],w[62],c[53],p[13],c[54]);
fulladd fa48(c[47],w[63],c[54],p[14],p[15]);
endmodule
module halfadd(a,b,sum,carry);
input a,b;
output sum,carry;
assign sum=a^b;
assign carry=a&b;
endmodule
module fulladd(a,b,c,sum,carry);
input a,b,c;
output sum,carry;
assign sum=a^b^c;
assign carry=(a&b)|(a&c)|(b&c);
endmodule
